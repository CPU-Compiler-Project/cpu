----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 09.05.2022 14:58:50
-- Design Name: 
-- Module Name: InstructionMemory - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity InstructionMemory is
    Port ( ADDR : in STD_LOGIC_VECTOR (7 downto 0);
           CLK : in STD_LOGIC;
           OUTPUT : out STD_LOGIC_VECTOR (31 downto 0));
end InstructionMemory;

architecture Behavioral of InstructionMemory is

type tabType is array(63 downto 0) of STD_LOGIC_VECTOR (31 downto 0);

signal instructionMem: tabType := ( -- THIS IS THE ROM : IT SHOULD CONTAINS THE CONTENT OF THE ASM FILE GENERATED BY OUR COMPILER
    X"00000004", -- @63 => AFC 0x1 (example)
    X"00000001", --
    X"00000002", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000000", --
    X"00000003" -- @0 => AFC 0x1 (example)
);

begin
    process(CLK) is
    begin
        if rising_edge(CLK) then
            OUTPUT <= instructionMem(to_integer(unsigned(ADDR)));
        end if;
    end process;

end Behavioral;
