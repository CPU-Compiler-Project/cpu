----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 09.05.2022 14:58:50
-- Design Name: 
-- Module Name: InstructionMemory - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity InstructionMemory is
    Port ( ADDR : in STD_LOGIC_VECTOR (7 downto 0);
           CLK : in STD_LOGIC;
           OUTPUT : out STD_LOGIC_VECTOR (31 downto 0));
end InstructionMemory;

architecture Behavioral of InstructionMemory is

type tabType is array(255 downto 0) of STD_LOGIC_VECTOR (31 downto 0);

signal instructionMem: tabType := ( -- THIS IS THE ROM : IT SHOULD CONTAINS THE CONTENT OF THE ASM FILE GENERATED BY OUR COMPILER
  X"00000000" -- @0xff
, X"00000000" -- @0xfe
, X"00000000" -- @0xfd
, X"00000000" -- @0xfc
, X"00000000" -- @0xfb
, X"00000000" -- @0xfa
, X"00000000" -- @0xf9
, X"00000000" -- @0xf8
, X"00000000" -- @0xf7
, X"00000000" -- @0xf6
, X"00000000" -- @0xf5
, X"00000000" -- @0xf4
, X"00000000" -- @0xf3
, X"00000000" -- @0xf2
, X"00000000" -- @0xf1
, X"00000000" -- @0xf0
, X"00000000" -- @0xef
, X"00000000" -- @0xee
, X"00000000" -- @0xed
, X"00000000" -- @0xec
, X"00000000" -- @0xeb
, X"00000000" -- @0xea
, X"00000000" -- @0xe9
, X"00000000" -- @0xe8
, X"00000000" -- @0xe7
, X"00000000" -- @0xe6
, X"00000000" -- @0xe5
, X"00000000" -- @0xe4
, X"00000000" -- @0xe3
, X"00000000" -- @0xe2
, X"00000000" -- @0xe1
, X"00000000" -- @0xe0
, X"00000000" -- @0xdf
, X"00000000" -- @0xde
, X"00000000" -- @0xdd
, X"00000000" -- @0xdc
, X"00000000" -- @0xdb
, X"00000000" -- @0xda
, X"00000000" -- @0xd9
, X"00000000" -- @0xd8
, X"00000000" -- @0xd7
, X"00000000" -- @0xd6
, X"00000000" -- @0xd5
, X"00000000" -- @0xd4
, X"00000000" -- @0xd3
, X"00000000" -- @0xd2
, X"00000000" -- @0xd1
, X"00000000" -- @0xd0
, X"00000000" -- @0xcf
, X"00000000" -- @0xce
, X"00000000" -- @0xcd
, X"00000000" -- @0xcc
, X"00000000" -- @0xcb
, X"00000000" -- @0xca
, X"00000000" -- @0xc9
, X"00000000" -- @0xc8
, X"00000000" -- @0xc7
, X"00000000" -- @0xc6
, X"00000000" -- @0xc5
, X"00000000" -- @0xc4
, X"00000000" -- @0xc3
, X"00000000" -- @0xc2
, X"00000000" -- @0xc1
, X"00000000" -- @0xc0
, X"00000000" -- @0xbf
, X"00000000" -- @0xbe
, X"00000000" -- @0xbd
, X"00000000" -- @0xbc
, X"00000000" -- @0xbb
, X"00000000" -- @0xba
, X"00000000" -- @0xb9
, X"00000000" -- @0xb8
, X"00000000" -- @0xb7
, X"00000000" -- @0xb6
, X"00000000" -- @0xb5
, X"00000000" -- @0xb4
, X"00000000" -- @0xb3
, X"00000000" -- @0xb2
, X"00000000" -- @0xb1
, X"00000000" -- @0xb0
, X"00000000" -- @0xaf
, X"00000000" -- @0xae
, X"00000000" -- @0xad
, X"00000000" -- @0xac
, X"00000000" -- @0xab
, X"00000000" -- @0xaa
, X"00000000" -- @0xa9
, X"00000000" -- @0xa8
, X"00000000" -- @0xa7
, X"00000000" -- @0xa6
, X"00000000" -- @0xa5
, X"00000000" -- @0xa4
, X"00000000" -- @0xa3
, X"00000000" -- @0xa2
, X"00000000" -- @0xa1
, X"00000000" -- @0xa0
, X"00000000" -- @0x9f
, X"00000000" -- @0x9e
, X"00000000" -- @0x9d
, X"00000000" -- @0x9c
, X"00000000" -- @0x9b
, X"00000000" -- @0x9a
, X"00000000" -- @0x99
, X"00000000" -- @0x98
, X"00000000" -- @0x97
, X"00000000" -- @0x96
, X"00000000" -- @0x95
, X"00000000" -- @0x94
, X"00000000" -- @0x93
, X"00000000" -- @0x92
, X"00000000" -- @0x91
, X"00000000" -- @0x90
, X"00000000" -- @0x8f
, X"00000000" -- @0x8e
, X"00000000" -- @0x8d
, X"00000000" -- @0x8c
, X"00000000" -- @0x8b
, X"00000000" -- @0x8a
, X"00000000" -- @0x89
, X"00000000" -- @0x88
, X"00000000" -- @0x87
, X"00000000" -- @0x86
, X"00000000" -- @0x85
, X"00000000" -- @0x84
, X"00000000" -- @0x83
, X"00000000" -- @0x82
, X"00000000" -- @0x81
, X"00000000" -- @0x80
, X"00000000" -- @0x7f
, X"00000000" -- @0x7e
, X"00000000" -- @0x7d
, X"00000000" -- @0x7c
, X"00000000" -- @0x7b
, X"00000000" -- @0x7a
, X"00000000" -- @0x79
, X"00000000" -- @0x78
, X"00000000" -- @0x77
, X"00000000" -- @0x76
, X"00000000" -- @0x75
, X"00000000" -- @0x74
, X"00000000" -- @0x73
, X"00000000" -- @0x72
, X"00000000" -- @0x71
, X"00000000" -- @0x70
, X"00000000" -- @0x6f
, X"00000000" -- @0x6e
, X"00000000" -- @0x6d
, X"00000000" -- @0x6c
, X"00000000" -- @0x6b
, X"00000000" -- @0x6a
, X"00000000" -- @0x69
, X"00000000" -- @0x68
, X"00000000" -- @0x67
, X"00000000" -- @0x66
, X"00000000" -- @0x65
, X"00000000" -- @0x64
, X"00000000" -- @0x63
, X"00000000" -- @0x62
, X"00000000" -- @0x61
, X"00000000" -- @0x60
, X"00000000" -- @0x5f
, X"00000000" -- @0x5e
, X"00000000" -- @0x5d
, X"00000000" -- @0x5c
, X"00000000" -- @0x5b
, X"00000000" -- @0x5a
, X"00000000" -- @0x59
, X"00000000" -- @0x58
, X"00000000" -- @0x57
, X"00000000" -- @0x56
, X"00000000" -- @0x55
, X"00000000" -- @0x54
, X"05121300" -- @0x53 => COP 0x12 0x13
, X"06130500" -- @0x52 => AFC 0x13 5
, X"06120000" -- @0x51 => AFC 0x12 0
, X"050a1200" -- @0x50 => COP 0x0a 0x12
, X"06120500" -- @0x4f => AFC 0x12 5
, X"06110000" -- @0x4e => AFC 0x11 0
, X"05101100" -- @0x4d => COP 0x10 0x11
, X"06110400" -- @0x4c => AFC 0x11 4
, X"06100000" -- @0x4b => AFC 0x10 0
, X"060f0000" -- @0x4a => AFC 0x0f 0
, X"090b0000" -- @0x49 => JMP 0x0b
, X"090d0000" -- @0x48 => JMP 0x0d
, X"090e0000" -- @0x47 => JMP 0x0e
, X"05010f00" -- @0x46 => COP 0x01 0x0f
, X"060f0000" -- @0x45 => AFC 0x0f 0
, X"0a480000" -- @0x44 => JMPF 0x48
, X"050e0100" -- @0x43 => COP 0x0e 0x01
, X"05000e00" -- @0x42 => COP 0x00 0x0e
, X"060e0000" -- @0x41 => AFC 0x0e 0
, X"0a490000" -- @0x40 => JMPF 0x49
, X"050d0000" -- @0x3f => COP 0x0d 0x00
, X"05000d00" -- @0x3e => COP 0x00 0x0d
, X"020d0d0e" -- @0x3d => MUL 0x0d 0x0d 0x0e
, X"050e0200" -- @0x3c => COP 0x0e 0x02
, X"050d0000" -- @0x3b => COP 0x0d 0x00
, X"0a3f0000" -- @0x3a => JMPF 0x3f
, X"050c0000" -- @0x39 => COP 0x0c 0x00
, X"05020c00" -- @0x38 => COP 0x02 0x0c
, X"060c0000" -- @0x37 => AFC 0x0c 0
, X"0a4a0000" -- @0x36 => JMPF 0x4a
, X"020b0b0c" -- @0x35 => MUL 0x0b 0x0b 0x0c
, X"060c0200" -- @0x34 => AFC 0x0c 2
, X"050b0200" -- @0x33 => COP 0x0b 0x02
, X"060a0000" -- @0x32 => AFC 0x0a 0
, X"09090000" -- @0x31 => JMP 0x09
, X"05000a00" -- @0x30 => COP 0x00 0x0a
, X"060a0000" -- @0x2f => AFC 0x0a 0
, X"0a320000" -- @0x2e => JMPF 0x32
, X"05090000" -- @0x2d => COP 0x09 0x00
, X"0a320000" -- @0x2c => JMPF 0x32
, X"05000900" -- @0x2b => COP 0x00 0x09
, X"0109090a" -- @0x2a => ADD 0x09 0x09 0x0a
, X"060a0200" -- @0x29 => AFC 0x0a 2
, X"05090000" -- @0x28 => COP 0x09 0x00
, X"0a2d0000" -- @0x27 => JMPF 0x2d
, X"01080809" -- @0x26 => ADD 0x08 0x08 0x09
, X"05090000" -- @0x25 => COP 0x09 0x00
, X"05080200" -- @0x24 => COP 0x08 0x02
, X"0a320000" -- @0x23 => JMPF 0x32
, X"06070000" -- @0x22 => AFC 0x07 0
, X"0a240000" -- @0x21 => JMPF 0x24
, X"06060000" -- @0x20 => AFC 0x06 0
, X"0a320000" -- @0x1f => JMPF 0x32
, X"06050000" -- @0x1e => AFC 0x05 0
, X"0a200000" -- @0x1d => JMPF 0x20
, X"05040100" -- @0x1c => COP 0x04 0x01
, X"05010400" -- @0x1b => COP 0x01 0x04
, X"06040000" -- @0x1a => AFC 0x04 0
, X"0a1c0000" -- @0x19 => JMPF 0x1c
, X"05010400" -- @0x18 => COP 0x01 0x04
, X"06040100" -- @0x17 => AFC 0x04 1
, X"0a1a0000" -- @0x16 => JMPF 0x1a
, X"02030304" -- @0x15 => MUL 0x03 0x03 0x04
, X"06040000" -- @0x14 => AFC 0x04 0
, X"06030100" -- @0x13 => AFC 0x03 1
, X"05000300" -- @0x12 => COP 0x00 0x03
, X"03030304" -- @0x11 => SOU 0x03 0x03 0x04
, X"06040500" -- @0x10 => AFC 0x04 5
, X"01030304" -- @0x0f => ADD 0x03 0x03 0x04
, X"04040405" -- @0x0e => DIV 0x04 0x04 0x05
, X"06050700" -- @0x0d => AFC 0x05 7
, X"02040405" -- @0x0c => MUL 0x04 0x04 0x05
, X"06050800" -- @0x0b => AFC 0x05 8
, X"06040900" -- @0x0a => AFC 0x04 9
, X"06030500" -- @0x09 => AFC 0x03 5
, X"05020300" -- @0x08 => COP 0x02 0x03
, X"06030500" -- @0x07 => AFC 0x03 5
, X"05020300" -- @0x06 => COP 0x02 0x03
, X"06035a00" -- @0x05 => AFC 0x03 90
, X"06020000" -- @0x04 => AFC 0x02 0
, X"06010000" -- @0x03 => AFC 0x01 0
, X"05000100" -- @0x02 => COP 0x00 0x01
, X"06010100" -- @0x01 => AFC 0x01 1
, X"06000000" -- @0x00 => AFC 0x00 0
);

begin
    process(CLK) is
    begin
        if rising_edge(CLK) then
            OUTPUT <= instructionMem(to_integer(unsigned(ADDR)));
        end if;
    end process;

end Behavioral;
