----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 09.05.2022 14:58:50
-- Design Name: 
-- Module Name: InstructionMemory - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity InstructionMemory is
    Port ( ADDR : in STD_LOGIC_VECTOR (7 downto 0);
           CLK : in STD_LOGIC;
           OUTPUT : out STD_LOGIC_VECTOR (31 downto 0));
end InstructionMemory;

architecture Behavioral of InstructionMemory is

type tabType is array(255 downto 0) of STD_LOGIC_VECTOR (31 downto 0);

signal instructionMem: tabType := ( -- THIS IS THE ROM : IT SHOULD CONTAINS THE CONTENT OF THE ASM FILE GENERATED BY OUR COMPILER
  X"00000000" -- @0xff
, X"00000000" -- @0xfe
, X"00000000" -- @0xfd
, X"00000000" -- @0xfc
, X"00000000" -- @0xfb
, X"00000000" -- @0xfa
, X"00000000" -- @0xf9
, X"00000000" -- @0xf8
, X"00000000" -- @0xf7
, X"00000000" -- @0xf6
, X"00000000" -- @0xf5
, X"00000000" -- @0xf4
, X"00000000" -- @0xf3
, X"00000000" -- @0xf2
, X"00000000" -- @0xf1
, X"00000000" -- @0xf0
, X"00000000" -- @0xef
, X"00000000" -- @0xee
, X"00000000" -- @0xed
, X"00000000" -- @0xec
, X"00000000" -- @0xeb
, X"00000000" -- @0xea
, X"00000000" -- @0xe9
, X"00000000" -- @0xe8
, X"00000000" -- @0xe7
, X"00000000" -- @0xe6
, X"00000000" -- @0xe5
, X"00000000" -- @0xe4
, X"00000000" -- @0xe3
, X"00000000" -- @0xe2
, X"00000000" -- @0xe1
, X"00000000" -- @0xe0
, X"00000000" -- @0xdf
, X"00000000" -- @0xde
, X"00000000" -- @0xdd
, X"00000000" -- @0xdc
, X"00000000" -- @0xdb
, X"00000000" -- @0xda
, X"00000000" -- @0xd9
, X"00000000" -- @0xd8
, X"00000000" -- @0xd7
, X"00000000" -- @0xd6
, X"00000000" -- @0xd5
, X"00000000" -- @0xd4
, X"00000000" -- @0xd3
, X"00000000" -- @0xd2
, X"00000000" -- @0xd1
, X"00000000" -- @0xd0
, X"00000000" -- @0xcf
, X"00000000" -- @0xce
, X"00000000" -- @0xcd
, X"00000000" -- @0xcc
, X"00000000" -- @0xcb
, X"00000000" -- @0xca
, X"00000000" -- @0xc9
, X"00000000" -- @0xc8
, X"00000000" -- @0xc7
, X"00000000" -- @0xc6
, X"00000000" -- @0xc5
, X"00000000" -- @0xc4
, X"00000000" -- @0xc3
, X"00000000" -- @0xc2
, X"00000000" -- @0xc1
, X"00000000" -- @0xc0
, X"00000000" -- @0xbf
, X"00000000" -- @0xbe
, X"00000000" -- @0xbd
, X"00000000" -- @0xbc
, X"00000000" -- @0xbb
, X"00000000" -- @0xba
, X"00000000" -- @0xb9
, X"00000000" -- @0xb8
, X"00000000" -- @0xb7
, X"00000000" -- @0xb6
, X"00000000" -- @0xb5
, X"00000000" -- @0xb4
, X"00000000" -- @0xb3
, X"00000000" -- @0xb2
, X"00000000" -- @0xb1
, X"00000000" -- @0xb0
, X"00000000" -- @0xaf
, X"00000000" -- @0xae
, X"00000000" -- @0xad
, X"00000000" -- @0xac
, X"00000000" -- @0xab
, X"00000000" -- @0xaa
, X"00000000" -- @0xa9
, X"00000000" -- @0xa8
, X"00000000" -- @0xa7
, X"00000000" -- @0xa6
, X"00000000" -- @0xa5
, X"00000000" -- @0xa4
, X"00000000" -- @0xa3
, X"00000000" -- @0xa2
, X"00000000" -- @0xa1
, X"00000000" -- @0xa0
, X"00000000" -- @0x9f
, X"00000000" -- @0x9e
, X"00000000" -- @0x9d
, X"00000000" -- @0x9c
, X"00000000" -- @0x9b
, X"00000000" -- @0x9a
, X"00000000" -- @0x99
, X"00000000" -- @0x98
, X"00000000" -- @0x97
, X"00000000" -- @0x96
, X"00000000" -- @0x95
, X"00000000" -- @0x94
, X"00000000" -- @0x93
, X"00000000" -- @0x92
, X"00000000" -- @0x91
, X"00000000" -- @0x90
, X"00000000" -- @0x8f
, X"00000000" -- @0x8e
, X"00000000" -- @0x8d
, X"00000000" -- @0x8c
, X"00000000" -- @0x8b
, X"00000000" -- @0x8a
, X"00000000" -- @0x89
, X"00000000" -- @0x88
, X"00000000" -- @0x87
, X"00000000" -- @0x86
, X"00000000" -- @0x85
, X"00000000" -- @0x84
, X"00000000" -- @0x83
, X"00000000" -- @0x82
, X"00000000" -- @0x81
, X"00000000" -- @0x80
, X"00000000" -- @0x7f
, X"00000000" -- @0x7e
, X"00000000" -- @0x7d
, X"00000000" -- @0x7c
, X"00000000" -- @0x7b
, X"00000000" -- @0x7a
, X"00000000" -- @0x79
, X"00000000" -- @0x78
, X"00000000" -- @0x77
, X"00000000" -- @0x76
, X"00000000" -- @0x75
, X"00000000" -- @0x74
, X"00000000" -- @0x73
, X"00000000" -- @0x72
, X"00000000" -- @0x71
, X"00000000" -- @0x70
, X"00000000" -- @0x6f
, X"00000000" -- @0x6e
, X"00000000" -- @0x6d
, X"00000000" -- @0x6c
, X"00000000" -- @0x6b
, X"00000000" -- @0x6a
, X"00000000" -- @0x69
, X"00000000" -- @0x68
, X"00000000" -- @0x67
, X"00000000" -- @0x66
, X"00000000" -- @0x65
, X"00000000" -- @0x64
, X"00000000" -- @0x63
, X"00000000" -- @0x62
, X"00000000" -- @0x61
, X"00000000" -- @0x60
, X"00000000" -- @0x5f
, X"00000000" -- @0x5e
, X"00000000" -- @0x5d
, X"00000000" -- @0x5c
, X"00000000" -- @0x5b
, X"00000000" -- @0x5a
, X"00000000" -- @0x59
, X"00000000" -- @0x58
, X"00000000" -- @0x57
, X"00000000" -- @0x56
, X"00000000" -- @0x55
, X"00000000" -- @0x54
, X"00000000" -- @0x53
, X"00000000" -- @0x52
, X"00000000" -- @0x51
, X"00000000" -- @0x50
, X"00000000" -- @0x4f
, X"00000000" -- @0x4e
, X"00000000" -- @0x4d
, X"00000000" -- @0x4c
, X"00000000" -- @0x4b
, X"00000000" -- @0x4a
, X"00000000" -- @0x49
, X"00000000" -- @0x48
, X"00000000" -- @0x47
, X"00000000" -- @0x46
, X"00000000" -- @0x45
, X"00000000" -- @0x44
, X"00000000" -- @0x43
, X"00000000" -- @0x42
, X"00000000" -- @0x41
, X"00000000" -- @0x40
, X"00000000" -- @0x3f
, X"00000000" -- @0x3e
, X"00000000" -- @0x3d
, X"00000000" -- @0x3c
, X"00000000" -- @0x3b
, X"00000000" -- @0x3a
, X"00000000" -- @0x39
, X"00000000" -- @0x38
, X"00000000" -- @0x37
, X"00000000" -- @0x36
, X"00000000" -- @0x35
, X"00000000" -- @0x34
, X"00000000" -- @0x33
, X"00000000" -- @0x32
, X"00000000" -- @0x31
, X"00000000" -- @0x30
, X"00000000" -- @0x2f
, X"00000000" -- @0x2e
, X"00000000" -- @0x2d
, X"00000000" -- @0x2c
, X"00000000" -- @0x2b
, X"00000000" -- @0x2a
, X"00000000" -- @0x29
, X"00000000" -- @0x28
, X"05070800" -- @0x27 => COP 0x07 0x08
, X"06080500" -- @0x26 => AFC 0x08 5
, X"06070000" -- @0x25 => AFC 0x07 0
, X"05030700" -- @0x24 => COP 0x03 0x07
, X"06070500" -- @0x23 => AFC 0x07 5
, X"06060000" -- @0x22 => AFC 0x06 0
, X"05050600" -- @0x21 => COP 0x05 0x06
, X"06060400" -- @0x20 => AFC 0x06 4
, X"06050000" -- @0x1f => AFC 0x05 0
, X"06040000" -- @0x1e => AFC 0x04 0
, X"05000400" -- @0x1d => COP 0x00 0x04
, X"02040405" -- @0x1c => MUL 0x04 0x04 0x05
, X"05050200" -- @0x1b => COP 0x05 0x02
, X"05040000" -- @0x1a => COP 0x04 0x00
, X"06030000" -- @0x19 => AFC 0x03 0
, X"05010300" -- @0x18 => COP 0x01 0x03
, X"01030304" -- @0x17 => ADD 0x03 0x03 0x04
, X"05040000" -- @0x16 => COP 0x04 0x00
, X"05030200" -- @0x15 => COP 0x03 0x02
, X"05010300" -- @0x14 => COP 0x01 0x03
, X"02030304" -- @0x13 => MUL 0x03 0x03 0x04
, X"06040000" -- @0x12 => AFC 0x04 0
, X"06030100" -- @0x11 => AFC 0x03 1
, X"05000300" -- @0x10 => COP 0x00 0x03
, X"03030304" -- @0x0f => SOU 0x03 0x03 0x04
, X"06040500" -- @0x0e => AFC 0x04 5
, X"01030304" -- @0x0d => ADD 0x03 0x03 0x04
, X"02040405" -- @0x0c => MUL 0x04 0x04 0x05
, X"06050800" -- @0x0b => AFC 0x05 8
, X"06040900" -- @0x0a => AFC 0x04 9
, X"06030500" -- @0x09 => AFC 0x03 5
, X"05020300" -- @0x08 => COP 0x02 0x03
, X"06030500" -- @0x07 => AFC 0x03 5
, X"05020300" -- @0x06 => COP 0x02 0x03
, X"06035a00" -- @0x05 => AFC 0x03 90
, X"06020000" -- @0x04 => AFC 0x02 0
, X"06010000" -- @0x03 => AFC 0x01 0
, X"05000100" -- @0x02 => COP 0x00 0x01
, X"06010100" -- @0x01 => AFC 0x01 1
, X"06000000" -- @0x00 => AFC 0x00 0
);

begin
    process(CLK) is
    begin
        if rising_edge(CLK) then
            OUTPUT <= instructionMem(to_integer(unsigned(ADDR)));
        end if;
    end process;

end Behavioral;
